bind v_bb_model v_bb_model_checker c0 (
    .CLK(CLK),
    .RST(RST),
    .REQ(REQ),
    .ACK(ACK),
    .OPCH(OPCH),
    .DONE(DONE),
    .ERR(ERR),
    .OPS(OPS),
    .TEST(TEST),
    .AB(AB),
    .BC(BC),
    .CD(CD),
    .BUSY(BUSY),
    .DATA(DATA),
    .STALL(STALL)
);

