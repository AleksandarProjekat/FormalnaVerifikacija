bind sv_model sv_model_checker c0 (
    .clk(clk),
    .rst(rst),
    .x(x),
    .y(y)

);

