bind black_box black_box_checker c0 (
    .clk(clk), .reset(reset),
    .a1(a1), .a2(a2), .a3(a3),
    .count_a(count_a), 
    .b(b),
    .c1(c1), .c2(c2), .c3(c3), .c4(c4),
    .a5(a5), .a6(a6),
    .b1(b1), .b2(b2), .b3(b3), .b4(b4)
);

